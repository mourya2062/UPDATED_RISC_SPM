`timescale 1ns / 1ps

module test_RISC_SPM ();
  reg rst;
  wire clk;
  parameter word_size = 8;
  reg [8:0] k;

  Clock_Unit M1 (clk);
  RISC_SPM M2 (clk, rst);

 initial #3500 $finish;
 
// Initialize Memory

initial begin
  #2 rst = 0; for (k=0;k<=255;k=k+1)M2.M2_SRAM.memory[k] = 0; #10 rst = 1;
end

initial begin
 

 #5
// opcode_src_dest
 M2.M2_SRAM.memory[0] = 8'b0000_00_00;		// NOP
 M2.M2_SRAM.memory[1] = 8'b0101_00_10;		// Read 130 to R2
 M2.M2_SRAM.memory[2] = 130;
 M2.M2_SRAM.memory[3] = 8'b0101_00_11;		// Read 131 to R3
 M2.M2_SRAM.memory[4] = 131;

 M2.M2_SRAM.memory[5] = 8'b1010_10_11;		// Multiply R2 and R3 and load R2 with Product_LSB and load R3 with product_MSB
 M2.M2_SRAM.memory[8] = 8'b0111_00_11;		// BR
 M2.M2_SRAM.memory[9] = 134;

// Load data
 M2.M2_SRAM.memory[130] = 5;
 M2.M2_SRAM.memory[131] = 6;
 M2.M2_SRAM.memory[134] = 139;
 M2.M2_SRAM.memory[139] = 8'b1111_00_00;		// HALT
 M2.M2_SRAM.memory[140] = 5;				//  Recycle
end 
//
endmodule 
